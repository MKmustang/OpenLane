`timescale 1ns / 1ps

module buffer (
    input wire in,
    output wire out
);

  assign out = in;

endmodule
